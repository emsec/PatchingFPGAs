module top(
    );

// top_earlgrey/u_rv_core_ibex/u_core/if_stage_i/gen_prefetch_buffer.prefetch_buffer_i/fifo_i/instr_addr_q_reg[%31..1%] : <- O
logic [30:0] instr_addr_i; // shifted by one bit to the right

// top_earlgrey/u_rv_core_ibex/u_core/if_stage_i/instr_out[%31..0%] : <- O
logic [31:0] instr_rdata_i;

// top_earlgrey/u_clkmgr/u_main_cg/i_cg/gen_xilinx.u_impl_xilinx/u_bufgce
logic clk_i;

logic [63:0] tinyla_probe;

assign tinyla_probe = {instr_addr_i, 1'b0, instr_rdata_i};

logic tinyla_trigger;

assign tinyla_trigger = (instr_addr_i == (32'h200003de >> 1)) ? 1'b1 : 1'b0;

typedef enum logic [1:0] {
STATE_RESET,
STATE_DO_SAMPLE,
STATE_IDLE
} tinyla_state_e;

logic [31:0] tinyla_doado;

logic [14:0] tinyla_buffer_read_addr;

logic [8:0] tinyla_buffer_write_addr;

logic bscan_drck;
logic bscan_reset;

logic tinyla_do_sample;

tinyla_state_e tinyla_state;
tinyla_state_e tinyla_state_next;

RAMB36E1 #(
// Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE" 
.RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
// Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
.SIM_COLLISION_CHECK("ALL"),
// DOA_REG, DOB_REG: Optional output register (0 or 1)
.DOA_REG(0),
.DOB_REG(0),
.EN_ECC_READ("FALSE"),                                                            // Enable ECC decoder,
                                                                                    // FALSE, TRUE
.EN_ECC_WRITE("FALSE"),                                                           // Enable ECC encoder,
                                                                                    // FALSE, TRUE
// INITP_00 to INITP_0F: Initial contents of the parity memory array
.INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
// INIT_00 to INIT_7F: Initial contents of the data memory array
.INIT_00(256'h8000000000000001800000000000000280000000000000038000000000000004),
.INIT_01(256'h8000000000000005800000000000000680000000000000078000000000000008),
.INIT_02(256'h8000000000000009800000000000000a800000000000000b800000000000000c),
.INIT_03(256'h800000000000000d800000000000000e800000000000000f8000000000000010),
.INIT_04(256'h8000000000000011800000000000001280000000000000138000000000000014),
.INIT_05(256'h8000000000000015800000000000001680000000000000178000000000000018),
.INIT_06(256'h8000000000000019800000000000001a800000000000001b800000000000001c),
.INIT_07(256'h800000000000001d800000000000001e800000000000001f8000000000000020),
.INIT_08(256'h8000000000000021800000000000002280000000000000238000000000000024),
.INIT_09(256'h8000000000000025800000000000002680000000000000278000000000000028),
.INIT_0A(256'h8000000000000029800000000000002a800000000000002b800000000000002c),
.INIT_0B(256'h800000000000002d800000000000002e800000000000002f8000000000000030),
.INIT_0C(256'h8000000000000031800000000000003280000000000000338000000000000034),
.INIT_0D(256'h8000000000000035800000000000003680000000000000378000000000000038),
.INIT_0E(256'h8000000000000039800000000000003a800000000000003b800000000000003c),
.INIT_0F(256'h800000000000003d800000000000003e800000000000003f8000000000000040),
.INIT_10(256'h8000000000000041800000000000004280000000000000438000000000000044),
.INIT_11(256'h8000000000000045800000000000004680000000000000478000000000000048),
.INIT_12(256'h8000000000000049800000000000004a800000000000004b800000000000004c),
.INIT_13(256'h800000000000004d800000000000004e800000000000004f8000000000000050),
.INIT_14(256'h8000000000000051800000000000005280000000000000538000000000000054),
.INIT_15(256'h8000000000000055800000000000005680000000000000578000000000000058),
.INIT_16(256'h8000000000000059800000000000005a800000000000005b800000000000005c),
.INIT_17(256'h800000000000005d800000000000005e800000000000005f8000000000000060),
.INIT_18(256'h8000000000000061800000000000006280000000000000638000000000000064),
.INIT_19(256'h8000000000000065800000000000006680000000000000678000000000000068),
.INIT_1A(256'h8000000000000069800000000000006a800000000000006b800000000000006c),
.INIT_1B(256'h800000000000006d800000000000006e800000000000006f8000000000000070),
.INIT_1C(256'h8000000000000071800000000000007280000000000000738000000000000074),
.INIT_1D(256'h8000000000000075800000000000007680000000000000778000000000000078),
.INIT_1E(256'h8000000000000079800000000000007a800000000000007b800000000000007c),
.INIT_1F(256'h800000000000007d800000000000007e800000000000007f8000000000000080),
.INIT_20(256'h8000000000000081800000000000008280000000000000838000000000000084),
.INIT_21(256'h8000000000000085800000000000008680000000000000878000000000000088),
.INIT_22(256'h8000000000000089800000000000008a800000000000008b800000000000008c),
.INIT_23(256'h800000000000008d800000000000008e800000000000008f8000000000000090),
.INIT_24(256'h8000000000000091800000000000009280000000000000938000000000000094),
.INIT_25(256'h8000000000000095800000000000009680000000000000978000000000000098),
.INIT_26(256'h8000000000000099800000000000009a800000000000009b800000000000009c),
.INIT_27(256'h800000000000009d800000000000009e800000000000009f80000000000000a0),
.INIT_28(256'h80000000000000a180000000000000a280000000000000a380000000000000a4),
.INIT_29(256'h80000000000000a580000000000000a680000000000000a780000000000000a8),
.INIT_2A(256'h80000000000000a980000000000000aa80000000000000ab80000000000000ac),
.INIT_2B(256'h80000000000000ad80000000000000ae80000000000000af80000000000000b0),
.INIT_2C(256'h80000000000000b180000000000000b280000000000000b380000000000000b4),
.INIT_2D(256'h80000000000000b580000000000000b680000000000000b780000000000000b8),
.INIT_2E(256'h80000000000000b980000000000000ba80000000000000bb80000000000000bc),
.INIT_2F(256'h80000000000000bd80000000000000be80000000000000bf80000000000000c0),
.INIT_30(256'h80000000000000c180000000000000c280000000000000c380000000000000c4),
.INIT_31(256'h80000000000000c580000000000000c680000000000000c780000000000000c8),
.INIT_32(256'h80000000000000c980000000000000ca80000000000000cb80000000000000cc),
.INIT_33(256'h80000000000000cd80000000000000ce80000000000000cf80000000000000d0),
.INIT_34(256'h80000000000000d180000000000000d280000000000000d380000000000000d4),
.INIT_35(256'h80000000000000d580000000000000d680000000000000d780000000000000d8),
.INIT_36(256'h80000000000000d980000000000000da80000000000000db80000000000000dc),
.INIT_37(256'h80000000000000dd80000000000000de80000000000000df80000000000000e0),
.INIT_38(256'h80000000000000e180000000000000e280000000000000e380000000000000e4),
.INIT_39(256'h80000000000000e580000000000000e680000000000000e780000000000000e8),
.INIT_3A(256'h80000000000000e980000000000000ea80000000000000eb80000000000000ec),
.INIT_3B(256'h80000000000000ed80000000000000ee80000000000000ef80000000000000f0),
.INIT_3C(256'h80000000000000f180000000000000f280000000000000f380000000000000f4),
.INIT_3D(256'h80000000000000f580000000000000f680000000000000f780000000000000f8),
.INIT_3E(256'h80000000000000f980000000000000fa80000000000000fb80000000000000fc),
.INIT_3F(256'h80000000000000fd80000000000000fe80000000000000ff8000000000000100),
.INIT_40(256'h8000000000000101800000000000010280000000000001038000000000000104),
.INIT_41(256'h8000000000000105800000000000010680000000000001078000000000000108),
.INIT_42(256'h8000000000000109800000000000010a800000000000010b800000000000010c),
.INIT_43(256'h800000000000010d800000000000010e800000000000010f8000000000000110),
.INIT_44(256'h8000000000000111800000000000011280000000000001138000000000000114),
.INIT_45(256'h8000000000000115800000000000011680000000000001178000000000000118),
.INIT_46(256'h8000000000000119800000000000011a800000000000011b800000000000011c),
.INIT_47(256'h800000000000011d800000000000011e800000000000011f8000000000000120),
.INIT_48(256'h8000000000000121800000000000012280000000000001238000000000000124),
.INIT_49(256'h8000000000000125800000000000012680000000000001278000000000000128),
.INIT_4A(256'h8000000000000129800000000000012a800000000000012b800000000000012c),
.INIT_4B(256'h800000000000012d800000000000012e800000000000012f8000000000000130),
.INIT_4C(256'h8000000000000131800000000000013280000000000001338000000000000134),
.INIT_4D(256'h8000000000000135800000000000013680000000000001378000000000000138),
.INIT_4E(256'h8000000000000139800000000000013a800000000000013b800000000000013c),
.INIT_4F(256'h800000000000013d800000000000013e800000000000013f8000000000000140),
.INIT_50(256'h8000000000000141800000000000014280000000000001438000000000000144),
.INIT_51(256'h8000000000000145800000000000014680000000000001478000000000000148),
.INIT_52(256'h8000000000000149800000000000014a800000000000014b800000000000014c),
.INIT_53(256'h800000000000014d800000000000014e800000000000014f8000000000000150),
.INIT_54(256'h8000000000000151800000000000015280000000000001538000000000000154),
.INIT_55(256'h8000000000000155800000000000015680000000000001578000000000000158),
.INIT_56(256'h8000000000000159800000000000015a800000000000015b800000000000015c),
.INIT_57(256'h800000000000015d800000000000015e800000000000015f8000000000000160),
.INIT_58(256'h8000000000000161800000000000016280000000000001638000000000000164),
.INIT_59(256'h8000000000000165800000000000016680000000000001678000000000000168),
.INIT_5A(256'h8000000000000169800000000000016a800000000000016b800000000000016c),
.INIT_5B(256'h800000000000016d800000000000016e800000000000016f8000000000000170),
.INIT_5C(256'h8000000000000171800000000000017280000000000001738000000000000174),
.INIT_5D(256'h8000000000000175800000000000017680000000000001778000000000000178),
.INIT_5E(256'h8000000000000179800000000000017a800000000000017b800000000000017c),
.INIT_5F(256'h800000000000017d800000000000017e800000000000017f8000000000000180),
.INIT_60(256'h8000000000000181800000000000018280000000000001838000000000000184),
.INIT_61(256'h8000000000000185800000000000018680000000000001878000000000000188),
.INIT_62(256'h8000000000000189800000000000018a800000000000018b800000000000018c),
.INIT_63(256'h800000000000018d800000000000018e800000000000018f8000000000000190),
.INIT_64(256'h8000000000000191800000000000019280000000000001938000000000000194),
.INIT_65(256'h8000000000000195800000000000019680000000000001978000000000000198),
.INIT_66(256'h8000000000000199800000000000019a800000000000019b800000000000019c),
.INIT_67(256'h800000000000019d800000000000019e800000000000019f80000000000001a0),
.INIT_68(256'h80000000000001a180000000000001a280000000000001a380000000000001a4),
.INIT_69(256'h80000000000001a580000000000001a680000000000001a780000000000001a8),
.INIT_6A(256'h80000000000001a980000000000001aa80000000000001ab80000000000001ac),
.INIT_6B(256'h80000000000001ad80000000000001ae80000000000001af80000000000001b0),
.INIT_6C(256'h80000000000001b180000000000001b280000000000001b380000000000001b4),
.INIT_6D(256'h80000000000001b580000000000001b680000000000001b780000000000001b8),
.INIT_6E(256'h80000000000001b980000000000001ba80000000000001bb80000000000001bc),
.INIT_6F(256'h80000000000001bd80000000000001be80000000000001bf80000000000001c0),
.INIT_70(256'h80000000000001c180000000000001c280000000000001c380000000000001c4),
.INIT_71(256'h80000000000001c580000000000001c680000000000001c780000000000001c8),
.INIT_72(256'h80000000000001c980000000000001ca80000000000001cb80000000000001cc),
.INIT_73(256'h80000000000001cd80000000000001ce80000000000001cf80000000000001d0),
.INIT_74(256'h80000000000001d180000000000001d280000000000001d380000000000001d4),
.INIT_75(256'h80000000000001d580000000000001d680000000000001d780000000000001d8),
.INIT_76(256'h80000000000001d980000000000001da80000000000001db80000000000001dc),
.INIT_77(256'h80000000000001dd80000000000001de80000000000001df80000000000001e0),
.INIT_78(256'h80000000000001e180000000000001e280000000000001e380000000000001e4),
.INIT_79(256'h80000000000001e580000000000001e680000000000001e780000000000001e8),
.INIT_7A(256'h80000000000001e980000000000001ea80000000000001eb80000000000001ec),
.INIT_7B(256'h80000000000001ed80000000000001ee80000000000001ef80000000000001f0),
.INIT_7C(256'h80000000000001f180000000000001f280000000000001f380000000000001f4),
.INIT_7D(256'h80000000000001f580000000000001f680000000000001f780000000000001f8),
.INIT_7E(256'h80000000000001f980000000000001fa80000000000001fb80000000000001fc),
.INIT_7F(256'h80000000000001fd80000000000001fe80000000000001ff8000000000000200),
// INIT_A, INIT_B: Initial values on output ports
.INIT_A(36'h000000000),
.INIT_B(36'h000000000),
// Initialization File: RAM initialization file
.INIT_FILE("NONE"),
// RAM Mode: "SDP" or "TDP" 
.RAM_MODE("SDP"),
// RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
.RAM_EXTENSION_A("NONE"),
.RAM_EXTENSION_B("NONE"),
// READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
.READ_WIDTH_A(1),                                                                 // 0-72
.READ_WIDTH_B(0),                                                                 // 0-36
.WRITE_WIDTH_A(0),                                                                // 0-36
.WRITE_WIDTH_B(72),                                                               // 0-72
// RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
.RSTREG_PRIORITY_A("RSTREG"),
.RSTREG_PRIORITY_B("RSTREG"),
// SRVAL_A, SRVAL_B: Set/reset value for output
.SRVAL_A(36'h000000000),
.SRVAL_B(36'h000000000),
// Simulation Device: Must be set to "7SERIES" for simulation behavior
.SIM_DEVICE("7SERIES"),
// WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
.WRITE_MODE_A("WRITE_FIRST"),
.WRITE_MODE_B("WRITE_FIRST")
)
tinyla_buffer (
// Cascade Signals: 1-bit (each) output: BRAM cascade ports (to create 64kx1)
.CASCADEOUTA(),                                   // 1-bit output: A port cascade
.CASCADEOUTB(),                                   // 1-bit output: B port cascade
// ECC Signals: 1-bit (each) output: Error Correction Circuitry ports
.DBITERR(),                                       // 1-bit output: Double bit error status
.ECCPARITY(),                                     // 8-bit output: Generated error correction parity
.RDADDRECC(),                                     // 9-bit output: ECC read address
.SBITERR(),                                       // 1-bit output: Single bit error status
// Port A Data: 32-bit (each) output: Port A data
.DOADO(tinyla_doado),                             // 32-bit output: A port data/LSB data
.DOPADOP(),                                       // 4-bit output: A port parity/LSB parity
// Port B Data: 32-bit (each) output: Port B data
.DOBDO(),                                         // 32-bit output: B port data/MSB data
.DOPBDOP(),                                       // 4-bit output: B port parity/MSB parity
// Cascade Signals: 1-bit (each) input: BRAM cascade ports (to create 64kx1)
.CASCADEINA(),                                    // 1-bit input: A port cascade
.CASCADEINB(),                                    // 1-bit input: B port cascade
// ECC Signals: 1-bit (each) input: Error Correction Circuitry ports
.INJECTDBITERR(),                                 // 1-bit input: Inject a double bit error
.INJECTSBITERR(),                                 // 1-bit input: Inject a single bit error
// Port A Address/Control Signals: 16-bit (each) input: Port A address and control signals (read port
// when RAM_MODE="SDP")
.ADDRARDADDR({1'b1, tinyla_buffer_read_addr}),    // 16-bit input: A port address/Read address
.CLKARDCLK(bscan_drck),                           // 1-bit input: A port clock/Read clock
.ENARDEN(1'b1),                                   // 1-bit input: A port enable/Read enable
.REGCEAREGCE(1'b0),                               // 1-bit input: A port register enable/Register enable
.RSTRAMARSTRAM(1'b0),                             // 1-bit input: A port set/reset
.RSTREGARSTREG(1'b0),                             // 1-bit input: A port register set/reset
.WEA(4'h0),                                       // 4-bit input: A port write enable
// Port A Data: 32-bit (each) input: Port A data
.DIADI(tinyla_probe[31:0]),                              // 32-bit input: A port data/LSB data
.DIPADIP(4'h0),                                   // 4-bit input: A port parity/LSB parity
// Port B Address/Control Signals: 16-bit (each) input: Port B address and control signals (write port
// when RAM_MODE="SDP")
.ADDRBWRADDR({1'b1, tinyla_buffer_write_addr, 6'h3f}),  // 16-bit input: B port address/Write address
.CLKBWRCLK(clk_i),                                  // 1-bit input: B port clock/Write clock
.ENBWREN(tinyla_do_sample),                       // 1-bit input: B port enable/Write enable
.REGCEB(1'b0),                                    // 1-bit input: B port register enable
.RSTRAMB(1'b0),                                   // 1-bit input: B port set/reset
.RSTREGB(1'b0),                                   // 1-bit input: B port register set/reset
.WEBWE(8'hff),                                    // 8-bit input: B port write enable/Write enable
// Port B Data: 32-bit (each) input: Port B data
.DIBDI(tinyla_probe[63:32]),                             // 32-bit input: B port data/MSB data
.DIPBDIP(4'h0)                                    // 4-bit input: B port parity/MSB parity
);

BSCANE2 #(
.JTAG_CHAIN(1)  // Value for USER command.
)
tinyla_jtag (
.CAPTURE(),                     // 1-bit output: CAPTURE output from TAP controller.
.DRCK(bscan_drck),              // 1-bit output: Gated TCK output. When SEL is asserted, DRCK toggles when CAPTURE or
                                // SHIFT are asserted.

.RESET(bscan_reset),            // 1-bit output: Reset output for TAP controller.
.RUNTEST(),                     // 1-bit output: Output asserted when TAP controller is in Run Test/Idle state.
.SEL(),                         // 1-bit output: USER instruction active output.
.SHIFT(),                       // 1-bit output: SHIFT output from TAP controller.
.TCK(),                         // 1-bit output: Test Clock output. Fabric connection to TAP Clock pin.
.TDI(),                         // 1-bit output: Test Data Input (TDI) output from TAP controller.
.TMS(),                         // 1-bit output: Test Mode Select output. Fabric connection to TAP.
.UPDATE(),                      // 1-bit output: UPDATE output from TAP controller
.TDO(tinyla_doado[0])           // 1-bit input: Test Data Output (TDO) input for USER function.
);

always_ff @(posedge bscan_drck or posedge bscan_reset) begin : tinyla_read_addr_cnt
if (bscan_reset) begin
    tinyla_buffer_read_addr <= 15'h0000;
end else begin
    tinyla_buffer_read_addr <= tinyla_buffer_read_addr + 1;
end
end

always_ff @(posedge clk_i or posedge bscan_reset) begin : tinyla_write_addr_cnt
if (bscan_reset) begin
    tinyla_buffer_write_addr <= 9'h000;
end else begin
    if (tinyla_do_sample) begin
    tinyla_buffer_write_addr <= tinyla_buffer_write_addr + 1;
    end
end
end

always_ff @(posedge clk_i or posedge bscan_reset) begin : tinyla_state_register
if (bscan_reset) begin
    tinyla_state <= STATE_RESET;
end else if ((tinyla_state == STATE_RESET && tinyla_trigger) || (tinyla_do_sample && tinyla_buffer_write_addr == 9'h1ff)) begin
    tinyla_state <= tinyla_state_next;
end
end

always_comb begin : tinyla_output_and_transition
unique case (tinyla_state)
    STATE_RESET:     tinyla_state_next = STATE_DO_SAMPLE;
    STATE_DO_SAMPLE: tinyla_state_next = STATE_IDLE;
    STATE_IDLE:      tinyla_state_next = STATE_IDLE;
    default:         tinyla_state_next = STATE_RESET;
endcase
end

assign tinyla_do_sample = (tinyla_state == STATE_DO_SAMPLE);

endmodule
